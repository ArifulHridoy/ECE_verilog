`timescale 1ns/10ps 
module tb; 
reg a, b; 
wire y; 
orgate uut (.a(a), .b(b), .y(y)); 
 
initial begin 
  $monitor("Time=%0t a=%b b=%b y=%b", $time, a, b, y); 
  $dumpfile("or.vcd"); 
  $dumpvars(0, tb); 
 
  a = 0; b = 0; 
  #10 a = 0; b = 1; 
  #10 a = 1; b = 0; 
  #10 a = 1; b = 1; 
  #10 $finish; 
end 
endmodule